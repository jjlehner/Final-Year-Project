module abc(
    input clk
);


endmodule : abc