module foo;

always_comb begin

end

endmodule : foo