module Pineapple (
    input logic jonah,
    output wire kathryn
);
logic fish;
endmodule