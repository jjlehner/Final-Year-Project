module foo;

initial begin
    block();
end

endmodule : foo