module foo;
    logic a;
    logic b;
endmodule : foo