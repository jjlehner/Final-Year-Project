module fish (
    input logic porty,
    output wire fishy
);

endmodule