module foo;
logic a;
endmodule : foo