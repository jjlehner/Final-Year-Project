module fish();

endmodule